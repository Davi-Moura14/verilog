module VERMELHO (

	input ckout,
	output VER

);

	assign VER = ckout; 
	
endmodule 